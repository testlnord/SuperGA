`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:20:13 04/01/2012 
// Design Name: 
// Module Name:    toAddr 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module toAddr(
// Global signals
    input wire ACLK,
//
    input wire [7:0] Xcoord,
    input wire [7:0] Ycoord,
	 output wire [7:0] Addr,
	 output wire Write
    );


endmodule
