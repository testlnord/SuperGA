`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:19:41 04/01/2012 
// Design Name: 
// Module Name:    toScreen 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module toScreen(
// Global signals
    input wire ACLK,
//
    input wire [7:0] Xcoord,
    input wire [7:0] Ycoord,
	 output wire [7:0] Xout,
	 output wire [7:0] Yout
    );


endmodule
